
--//32-bit CLA Behavioral Design//---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
-------------------------------------------------------------------------------------------------------------------------
entity CLA32_bh is
  port (A_32b: in std_logic_vector (31 downto 0);
        B_32b: in std_logic_vector (31 downto 0);
        C0_32b: in std_logic;
        S_32b: out std_logic_vector (31 downto 0);
	P_32b: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	G_32b: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
        C32_32b: out STD_LOGIC
        );
end CLA32_bh;
------------------------------------------------------------------------------------------------------------------------- 
architecture CLA32_behavioral of CLA32_bh is
-------------------------------------------------------------------------------------------------------------------------
--SIGNAL C4_32b,C8_32b, C12_32b,C16_32b: STD_LOGIC;
--SIGNAL C123_32b: STD_LOGIC_VECTOR (31 DOWNTO 0);
-------------------------------------------------------------------------------------------------------------------------
BEGIN
S_32b <= (A_32b + B_32b) + C0_32b;
end CLA32_behavioral;
-------------------------------------------------------------------------------------------------------------------------
